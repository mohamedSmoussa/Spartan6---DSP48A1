module DSP48A1 (A,B,C,D,BCIN,CARRYIN,M,P,CARRYOUT,CARRYOUTF,CLK,OPMODE,CEA,CEB,CEC,CECARRYIN,CED,CEM
                ,CEOPMODE,CEP,RSTA,RSTB,RSTC,RSTCARRYIN,RSTD,RSTM,RSTOPMODE,RSTP,BCOUT,PCIN,PCOUT);
parameter A0REG=0; parameter A1REG=1; parameter B0REG=0; parameter B1REG=1; parameter CREG=1;
parameter DREG=1; parameter MREG=1; parameter PREG=1;  parameter CAARYINREG=1; parameter CAARYOUTREG=1;
parameter OPMODEREG=1; parameter CARRYINSEL="OPMODE5"; parameter B_INPUT = "DIRECT"; parameter RSTTYPE = "SYNC" ;
input [17:0] A,B,D,BCIN;
input [47:0] C,PCIN;
input [7:0] OPMODE;
input CARRYIN,CLK,CEA,CEB,CEC,CECARRYIN,CED,CEM,CEOPMODE,CEP;
input RSTA,RSTB,RSTC,RSTCARRYIN,RSTD,RSTM,RSTOPMODE,RSTP;
output  [17:0] BCOUT ;
output [47:0]P,PCOUT;
output [35:0]M;
output  CARRYOUT,CARRYOUTF;
wire [17:0] MUXED_B,B0_S,A0_S,D_S,A1_S,PRE_OUT,B1_INPUT,B1_S;
wire [47:0] C_S,MUX_X_IN3,MUX_X_OUT,MUX_Z_OUT,POST_OUT,M_TO_MUX;
wire [7:0] OPMODE_S;
wire [35:0]MULT_OUT,M_S;
wire CARRYIN_S1,CIN,POST_COUT;
assign BCOUT=B1_S;
assign M=M_S;
assign PCOUT=P;
assign CARRYOUTF=CARRYOUT;
assign MUX_X_IN3={D_S[11:0],A1_S,B1_S};
assign M_TO_MUX={12'h000,M_S};
assign MUXED_B=(B_INPUT=="DIRECT")?B:(B_INPUT=="CASCADE")?BCIN:0;
assign CARRYIN_S1=(CARRYINSEL=="OPMODE5")?OPMODE_S[5]:(CARRYINSEL=="CARRYIN")?CARRYIN:0;
assign B1_INPUT=(OPMODE_S[4])?PRE_OUT:B0_S;
assign MULT_OUT=A1_S*B1_S;
assign PRE_OUT=(OPMODE_S[6])?D_S-B0_S:B0_S+D_S;
assign {POST_COUT,POST_OUT}=(OPMODE_S[7])? MUX_Z_OUT-(MUX_X_OUT+CIN):MUX_X_OUT+MUX_Z_OUT+CIN;
 MUX_REG_INPUT #(.WIDTH(8),.MODE(RSTTYPE)) OPMODE_SEL(OPMODE,OPMODEREG,OPMODE_S,CLK,RSTOPMODE,CEOPMODE);
 MUX_REG_INPUT #(.WIDTH(18),.MODE(RSTTYPE)) B0_SEL(MUXED_B,B0REG,B0_S,CLK,RSTB,CEB);
 MUX_REG_INPUT #(.WIDTH(18),.MODE(RSTTYPE)) A0_SEL(A,A0REG,A0_S,CLK,RSTA,CEA);
 MUX_REG_INPUT #(.WIDTH(18),.MODE(RSTTYPE)) A1_SEL(A0_S,A1REG,A1_S,CLK,RSTA,CEA);
 MUX_REG_INPUT #(.WIDTH(18),.MODE(RSTTYPE)) D_SEL(D,DREG,D_S,CLK,RSTD,CED);
 MUX_REG_INPUT #(.WIDTH(48),.MODE(RSTTYPE)) C_SEL(C,CREG,C_S,CLK,RSTC,CEC);
 MUX_REG_INPUT #(.WIDTH(18),.MODE(RSTTYPE)) B1_SEL(B1_INPUT,B1REG,B1_S,CLK,RSTB,CEB);
 MUX_REG_INPUT #(.WIDTH(36),.MODE(RSTTYPE)) M_SEL(MULT_OUT,MREG,M_S,CLK,RSTM,CEM);
 MUX4_1 #(.WIDTH(48)) MUX_X(M_TO_MUX,PCOUT,MUX_X_IN3,OPMODE_S[1:0],MUX_X_OUT);
 MUX4_1 #(.WIDTH(48)) MUX_Z(PCIN,PCOUT,C_S,OPMODE_S[3:2],MUX_Z_OUT);
 MUX_REG_INPUT #(.MODE(RSTTYPE)) CARRYIN_SEL(CARRYIN_S1,CAARYINREG,CIN,CLK,RSTCARRYIN,CECARRYIN);
 MUX_REG_INPUT #(.WIDTH(48),.MODE(RSTTYPE)) P_SEL(POST_OUT,PREG,P,CLK,RSTP,CEP);
 MUX_REG_INPUT #(.MODE(RSTTYPE)) CARRYOUT_SEL(POST_COUT,CAARYOUTREG,CARRYOUT,CLK,RSTCARRYIN,CECARRYIN);
endmodule //DSP48A1